module animate();